

module MMU #(
    parameter ADDR_WIDTH = 64
) (
    
)
    typedef logic[ADDR_WIDTH-1:0] addr_t;




endmodule