`ifndef __REG_STRUCT__
`define __REG_STRUCT__
package RegStruct;
    typedef struct {logic [63:0] regs[31:0];} RegPack;
endpackage
`endif
